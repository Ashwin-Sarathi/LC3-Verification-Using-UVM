//----------------------------------------------------------------------
// Created with uvmf_gen version 2023.4
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: 
// This file contains defines and typedefs to be compiled for use in
// the simulation running on the emulator when using Veloce.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
                                                                               

typedef bit enableWB_status_t;
typedef bit [2:0] psr_t;
typedef bit [15:0] VSR1_t;
typedef bit [15:0] VSR2_t;

// pragma uvmf custom additional begin
// pragma uvmf custom additional end

